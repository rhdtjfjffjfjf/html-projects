library IEEE
use IEEE.std_logic_1164.all;

Entity the_mux is port
(
	