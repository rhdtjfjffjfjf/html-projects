library IEEE;
use IEEE.std_logic_1164.all;

Entity my9bit is
end my9bit;

Architecture my9bita of my9bit is

component my8bit is port (
	   A: in std_logic_vector(7 downto 0);
		Y0: out std_logic_vector(7 downto 0);
		Y1: out std_logic_vector(7 downto 0);
		Y2: out Std_logic_vector(7 downto 0);
		Y3: out Std_logic_vector(7 downto 0);
		sel: in std_logic_vector(1 downto 0)
		);
end component;


signal sel1: std_logic_vector(1 downto 0);

Begin

DUT: my8bit port map(sel <= sel1);

sel1 <= "00", "01" after 50 ps, "10" after 100ps, "11" after 150ps;

end my9bita;







